library verilog;
use verilog.vl_types.all;
entity PrescalerTen_vlg_check_tst is
    port(
        clk_out         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end PrescalerTen_vlg_check_tst;
