library verilog;
use verilog.vl_types.all;
entity PrescalerSix_vlg_vec_tst is
end PrescalerSix_vlg_vec_tst;
