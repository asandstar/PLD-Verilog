library verilog;
use verilog.vl_types.all;
entity TimeCounter_vlg_vec_tst is
end TimeCounter_vlg_vec_tst;
