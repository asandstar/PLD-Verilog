library verilog;
use verilog.vl_types.all;
entity Washmachine_vlg_vec_tst is
end Washmachine_vlg_vec_tst;
