library verilog;
use verilog.vl_types.all;
entity WashmachineControl_vlg_vec_tst is
end WashmachineControl_vlg_vec_tst;
