library verilog;
use verilog.vl_types.all;
entity PrescalerTen_vlg_vec_tst is
end PrescalerTen_vlg_vec_tst;
