library verilog;
use verilog.vl_types.all;
entity SegDecode_vlg_vec_tst is
end SegDecode_vlg_vec_tst;
