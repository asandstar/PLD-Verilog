library verilog;
use verilog.vl_types.all;
entity DynamicScan_vlg_vec_tst is
end DynamicScan_vlg_vec_tst;
