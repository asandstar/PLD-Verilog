library verilog;
use verilog.vl_types.all;
entity PrescalerFour_vlg_vec_tst is
end PrescalerFour_vlg_vec_tst;
